library IEEE; 
 
use IEEE.std_logic_1164.all; 
--Additional standard or custom libraries go here 
 
package graphic_const is 
 	 
	
	constant TANK_WIDTH : natural := 80;
	constant TANK_HEIGHT  : natural := 60;
	constant BARREL_WIDTH : natural := 10;
	constant BARREL_HEIGHT : natural := 30;
 
 	--Other constants, types, subroutines, components go here 
 
end package graphic_const; 
 
package body graphic_const is 
 
--Subroutine declarations go here 
-- you will not have any need for it now, this package is only for defining -
-- some useful constants  
 
end package body graphic_const; 